module BCD10_4to2(
    input logic [3:0] b,
    output logic [7:0] p
    );
    always_comb
    case(b)
        //ʮ�������ֵ���ʾ
        4'b0000 : p = 8'b00000000;
        4'b0001 : p = 8'b00000001;
        4'b0010 : p = 8'b00000010;
        4'b0011 : p = 8'b00000011;
        4'b0100 : p = 8'b00000100;
        4'b0101 : p = 8'b00000101;
        4'b0110 : p = 8'b00000110;
        4'b0111 : p = 8'b00000111;
        4'b1000 : p = 8'b00001000;
        4'b1001 : p = 8'b00001001;
        4'b1010 : p = 8'b00010000;
        4'b1011 : p = 8'b00010001;
        4'b1100 : p = 8'b00010010;
        4'b1101 : p = 8'b00010011;
        4'b1110 : p = 8'b00010100;
        4'b1111 : p = 8'b00010101;
      endcase
endmodule
